    -- User Interface
    note_in <= note_next;
 
    process (CLK,RST) 
        variable state: integer range 0 to 100 := 0;
        variable del_cnt : integer range 0 to 1000000000 := 0;
        
        -- define an array of note values
        type note_array is array (natural range <>) of std_logic_vector(4 downto 0);
        constant song_notes : note_array := ("10001", "00000", "01100", "00000", "01010", "00000", "00101", "00000", "00101", "00000", "00101", "00000", "00101", "00000", "00101", "00000", "01010", "00000", "01010", "00000", "01010", "00000", "01010", "00000", "01010", "00000", "01000", "00000", "01010", "00000", "00110", "00000", "00110", "00000", "00110", "00000", "00110", "00000", "00110", "00000", "01010", "00000", "01010", "00000", "01010", "00000", "01010", "00000", "01010", "00000", "01100", "00000", "10001", "00000", "01000", "00000", "01000", "00000", "01000", "00000", "01000", "00000", "01000", "00000", "01000", "00000", "01000", "00000", "10001", "00000", "10001", "00000", "10001", "00000", "10011", "00000", "10011", "00000", "01100", "00000");
        -- define an array of delay values
        type delay_array is array (natural range <>) of integer;
        constant song_delays : delay_array := (32608695, 32608695, 32608695, 32608695, 16304347, 16304347, 16304347, 16304347, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 8152173, 16304347, 16304347, 16304347, 16304347, 16304347, 16304347, 97826086, 9782608);
    begin
        if (RST = '1') then
            state := 0;
            del_cnt := 0;
        elsif (CLK'event and CLK = '1') then
            if (del_cnt = 0 ) then
                -- iterate through the note and delay arrays
                note_next <= song_notes(state);
                del_cnt := song_delays(state);
                state := state + 1;
                
                -- reset the state to 0 when the end of the song is reached
                if (state = song_notes'length +1) then
                    state := 0;
                    del_cnt := 0;
                end if;
            else
                del_cnt := del_cnt - 1;
            end if;
        end if;
    end process;
    
end Behavioral;
